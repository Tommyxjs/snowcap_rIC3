module OneHotLatch #(
) (
input wire clk,
input wire [405:0] x,
output wire prop
);

    wire valid_input;
wire done;
reg [405:0] l;

    assign valid_input = (x != 0) && ((x & (x - 1)) == 0);
assign done = (l == 406'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111);
assign prop = done;

    always @(*) begin
assume(valid_input);
end

    always @(posedge clk) begin
l <= l | x;
end

    always @(*) begin
assume(!(x[15] && !(l[391] || l[383] || l[323])));
end

    always @(*) begin
assume(!(x[370] && !(l[293])));
end

    always @(*) begin
assume(!(x[293] && !(l[15])));
end

endmodule
