module OneHotLatch #()
(input wire clk,
input wire [2015:0] x,
output wire prop
);

    wire valid_input;
wire done;
reg [2015:0] l;
reg assume_failed;

    reg l2015_prev;
    reg l2000_prev;

    assign valid_input = (x != 0) && ((x & (x - 1)) == 0);
assign done = (l == 2016'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111);
assign prop = done;
wire assume_ok = !assume_failed;

    always @(*) begin
assume(valid_input);
end
always @(*) begin
assume(assume_ok);
end

    always @(posedge clk) begin
l <= l | x;
end

    always @(posedge clk) begin
if (valid_input && l[686] && !(l2015_prev || l2000_prev))
assume_failed <= 1;
        l2015_prev <= l[2015];
        l2000_prev <= l[2000];
    end

endmodule
